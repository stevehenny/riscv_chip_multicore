localparam RTYPEOP = 7'b0110011;
localparam ITYPEOP = 7'b0010011;
localparam ADDFUNCT3 = 3'b000;
localparam ADDFUNCT7 = 7'b0000000;
localparam SUBFUNCT3 = 3'b000;
localparam SUBFUNCT7 = 7'b0100000;
localparam ANDFUNCT3 = 3'b111;
localparam ANDFUNCT7 = 7'b0000000;
localparam ORFUNCT3 = 3'b110;
localparam ORFUNCT7 = 7'b0000000;
localparam XORFUNCT3 = 3'b100;
localparam XORFUNCT7 = 7'b0000000;
localparam SLLFUNCT3 = 3'b001;
localparam SLLFUNCT7 = 7'b0000000;
localparam SRLFUNCT3 = 3'b101;
localparam SRLFUNCT7 = 7'b0000000;
localparam SRAFUNCT3 = 3'b101;
localparam SRAFUNCT7 = 7'b0100000;
localparam SLTFUNCT3 = 3'b010;
localparam SLTFUNCT7 = 7'b0000000;
localparam SLTUFUNCT3 = 3'b011;
localparam SLTUFUNCT7 = 7'b0000000;
localparam MULFUNCT3 = 3'b000;
localparam MULFUNCT7 = 7'b0000001;
localparam DIVFUNCT7 = 7'b0000001;
localparam REMFUNCT7 = 7'b0000001;
